
module correction_lut_16(value, corrected); 

input [7:0] value; 
output [15:0] corrected; 
reg [15:0] corrected; 

always @(value) 

case (value) 
0: corrected=0;
1: corrected=3;
2: corrected=10;
3: corrected=22;
4: corrected=37;
5: corrected=55;
6: corrected=76;
7: corrected=101;
8: corrected=128;
9: corrected=159;
10: corrected=192;
11: corrected=228;
12: corrected=267;
13: corrected=308;
14: corrected=352;
15: corrected=399;
16: corrected=448;
17: corrected=500;
18: corrected=554;
19: corrected=611;
20: corrected=670;
21: corrected=732;
22: corrected=796;
23: corrected=862;
24: corrected=931;
25: corrected=1002;
26: corrected=1075;
27: corrected=1151;
28: corrected=1229;
29: corrected=1309;
30: corrected=1391;
31: corrected=1476;
32: corrected=1563;
33: corrected=1652;
34: corrected=1743;
35: corrected=1836;
36: corrected=1932;
37: corrected=2029;
38: corrected=2129;
39: corrected=2231;
40: corrected=2335;
41: corrected=2441;
42: corrected=2550;
43: corrected=2660;
44: corrected=2772;
45: corrected=2887;
46: corrected=3003;
47: corrected=3122;
48: corrected=3242;
49: corrected=3365;
50: corrected=3490;
51: corrected=3616;
52: corrected=3745;
53: corrected=3876;
54: corrected=4008;
55: corrected=4143;
56: corrected=4279;
57: corrected=4418;
58: corrected=4559;
59: corrected=4701;
60: corrected=4845;
61: corrected=4992;
62: corrected=5140;
63: corrected=5290;
64: corrected=5442;
65: corrected=5596;
66: corrected=5752;
67: corrected=5910;
68: corrected=6070;
69: corrected=6232;
70: corrected=6395;
71: corrected=6560;
72: corrected=6728;
73: corrected=6897;
74: corrected=7068;
75: corrected=7241;
76: corrected=7415;
77: corrected=7592;
78: corrected=7770;
79: corrected=7951;
80: corrected=8133;
81: corrected=8317;
82: corrected=8502;
83: corrected=8690;
84: corrected=8879;
85: corrected=9070;
86: corrected=9263;
87: corrected=9458;
88: corrected=9655;
89: corrected=9853;
90: corrected=10053;
91: corrected=10255;
92: corrected=10459;
93: corrected=10665;
94: corrected=10872;
95: corrected=11081;
96: corrected=11292;
97: corrected=11505;
98: corrected=11719;
99: corrected=11935;
100: corrected=12153;
101: corrected=12373;
102: corrected=12594;
103: corrected=12817;
104: corrected=13042;
105: corrected=13269;
106: corrected=13497;
107: corrected=13727;
108: corrected=13959;
109: corrected=14192;
110: corrected=14428;
111: corrected=14665;
112: corrected=14903;
113: corrected=15144;
114: corrected=15386;
115: corrected=15629;
116: corrected=15875;
117: corrected=16122;
118: corrected=16371;
119: corrected=16622;
120: corrected=16874;
121: corrected=17128;
122: corrected=17383;
123: corrected=17641;
124: corrected=17900;
125: corrected=18160;
126: corrected=18423;
127: corrected=18687;
128: corrected=18953;
129: corrected=19220;
130: corrected=19489;
131: corrected=19760;
132: corrected=20032;
133: corrected=20306;
134: corrected=20582;
135: corrected=20859;
136: corrected=21138;
137: corrected=21418;
138: corrected=21701;
139: corrected=21985;
140: corrected=22270;
141: corrected=22557;
142: corrected=22846;
143: corrected=23136;
144: corrected=23428;
145: corrected=23722;
146: corrected=24017;
147: corrected=24314;
148: corrected=24613;
149: corrected=24913;
150: corrected=25215;
151: corrected=25518;
152: corrected=25823;
153: corrected=26130;
154: corrected=26438;
155: corrected=26748;
156: corrected=27059;
157: corrected=27372;
158: corrected=27687;
159: corrected=28003;
160: corrected=28321;
161: corrected=28640;
162: corrected=28961;
163: corrected=29284;
164: corrected=29608;
165: corrected=29934;
166: corrected=30261;
167: corrected=30590;
168: corrected=30921;
169: corrected=31253;
170: corrected=31587;
171: corrected=31922;
172: corrected=32259;
173: corrected=32597;
174: corrected=32937;
175: corrected=33278;
176: corrected=33622;
177: corrected=33966;
178: corrected=34312;
179: corrected=34660;
180: corrected=35009;
181: corrected=35360;
182: corrected=35713;
183: corrected=36067;
184: corrected=36422;
185: corrected=36779;
186: corrected=37138;
187: corrected=37498;
188: corrected=37860;
189: corrected=38223;
190: corrected=38588;
191: corrected=38954;
192: corrected=39322;
193: corrected=39692;
194: corrected=40063;
195: corrected=40435;
196: corrected=40809;
197: corrected=41185;
198: corrected=41562;
199: corrected=41940;
200: corrected=42320;
201: corrected=42702;
202: corrected=43085;
203: corrected=43470;
204: corrected=43856;
205: corrected=44244;
206: corrected=44633;
207: corrected=45024;
208: corrected=45416;
209: corrected=45810;
210: corrected=46205;
211: corrected=46602;
212: corrected=47000;
213: corrected=47400;
214: corrected=47801;
215: corrected=48204;
216: corrected=48609;
217: corrected=49014;
218: corrected=49422;
219: corrected=49831;
220: corrected=50241;
221: corrected=50653;
222: corrected=51066;
223: corrected=51481;
224: corrected=51897;
225: corrected=52315;
226: corrected=52734;
227: corrected=53155;
228: corrected=53577;
229: corrected=54001;
230: corrected=54426;
231: corrected=54853;
232: corrected=55281;
233: corrected=55711;
234: corrected=56142;
235: corrected=56574;
236: corrected=57008;
237: corrected=57444;
238: corrected=57881;
239: corrected=58319;
240: corrected=58759;
241: corrected=59201;
242: corrected=59644;
243: corrected=60088;
244: corrected=60534;
245: corrected=60981;
246: corrected=61430;
247: corrected=61880;
248: corrected=62332;
249: corrected=62785;
250: corrected=63240;
251: corrected=63696;
252: corrected=64153;
253: corrected=64612;
254: corrected=65073;
255: corrected=65535;


endcase 

endmodule

