
module correction_lut_8(value, corrected); 

input [7:0] value; 
output [7:0] corrected; 
reg [7:0] corrected; 

always @(value) 

case (value) 
0: corrected=0;
1: corrected=0;
2: corrected=0;
3: corrected=0;
4: corrected=0;
5: corrected=0;
6: corrected=0;
7: corrected=0;
8: corrected=0;
9: corrected=0;
10: corrected=0;
11: corrected=0;
12: corrected=1;
13: corrected=1;
14: corrected=1;
15: corrected=1;
16: corrected=1;
17: corrected=1;
18: corrected=2;
19: corrected=2;
20: corrected=2;
21: corrected=2;
22: corrected=3;
23: corrected=3;
24: corrected=3;
25: corrected=3;
26: corrected=4;
27: corrected=4;
28: corrected=4;
29: corrected=5;
30: corrected=5;
31: corrected=5;
32: corrected=6;
33: corrected=6;
34: corrected=6;
35: corrected=7;
36: corrected=7;
37: corrected=7;
38: corrected=8;
39: corrected=8;
40: corrected=9;
41: corrected=9;
42: corrected=9;
43: corrected=10;
44: corrected=10;
45: corrected=11;
46: corrected=11;
47: corrected=12;
48: corrected=12;
49: corrected=13;
50: corrected=13;
51: corrected=14;
52: corrected=14;
53: corrected=15;
54: corrected=15;
55: corrected=16;
56: corrected=16;
57: corrected=17;
58: corrected=17;
59: corrected=18;
60: corrected=18;
61: corrected=19;
62: corrected=20;
63: corrected=20;
64: corrected=21;
65: corrected=21;
66: corrected=22;
67: corrected=22;
68: corrected=23;
69: corrected=24;
70: corrected=24;
71: corrected=25;
72: corrected=26;
73: corrected=26;
74: corrected=27;
75: corrected=28;
76: corrected=28;
77: corrected=29;
78: corrected=30;
79: corrected=30;
80: corrected=31;
81: corrected=32;
82: corrected=33;
83: corrected=33;
84: corrected=34;
85: corrected=35;
86: corrected=36;
87: corrected=36;
88: corrected=37;
89: corrected=38;
90: corrected=39;
91: corrected=39;
92: corrected=40;
93: corrected=41;
94: corrected=42;
95: corrected=43;
96: corrected=43;
97: corrected=44;
98: corrected=45;
99: corrected=46;
100: corrected=47;
101: corrected=48;
102: corrected=49;
103: corrected=49;
104: corrected=50;
105: corrected=51;
106: corrected=52;
107: corrected=53;
108: corrected=54;
109: corrected=55;
110: corrected=56;
111: corrected=57;
112: corrected=57;
113: corrected=58;
114: corrected=59;
115: corrected=60;
116: corrected=61;
117: corrected=62;
118: corrected=63;
119: corrected=64;
120: corrected=65;
121: corrected=66;
122: corrected=67;
123: corrected=68;
124: corrected=69;
125: corrected=70;
126: corrected=71;
127: corrected=72;
128: corrected=73;
129: corrected=74;
130: corrected=75;
131: corrected=76;
132: corrected=77;
133: corrected=79;
134: corrected=80;
135: corrected=81;
136: corrected=82;
137: corrected=83;
138: corrected=84;
139: corrected=85;
140: corrected=86;
141: corrected=87;
142: corrected=88;
143: corrected=90;
144: corrected=91;
145: corrected=92;
146: corrected=93;
147: corrected=94;
148: corrected=95;
149: corrected=96;
150: corrected=98;
151: corrected=99;
152: corrected=100;
153: corrected=101;
154: corrected=102;
155: corrected=104;
156: corrected=105;
157: corrected=106;
158: corrected=107;
159: corrected=108;
160: corrected=110;
161: corrected=111;
162: corrected=112;
163: corrected=113;
164: corrected=115;
165: corrected=116;
166: corrected=117;
167: corrected=119;
168: corrected=120;
169: corrected=121;
170: corrected=122;
171: corrected=124;
172: corrected=125;
173: corrected=126;
174: corrected=128;
175: corrected=129;
176: corrected=130;
177: corrected=132;
178: corrected=133;
179: corrected=134;
180: corrected=136;
181: corrected=137;
182: corrected=138;
183: corrected=140;
184: corrected=141;
185: corrected=143;
186: corrected=144;
187: corrected=145;
188: corrected=147;
189: corrected=148;
190: corrected=150;
191: corrected=151;
192: corrected=153;
193: corrected=154;
194: corrected=155;
195: corrected=157;
196: corrected=158;
197: corrected=160;
198: corrected=161;
199: corrected=163;
200: corrected=164;
201: corrected=166;
202: corrected=167;
203: corrected=169;
204: corrected=170;
205: corrected=172;
206: corrected=173;
207: corrected=175;
208: corrected=176;
209: corrected=178;
210: corrected=179;
211: corrected=181;
212: corrected=182;
213: corrected=184;
214: corrected=185;
215: corrected=187;
216: corrected=189;
217: corrected=190;
218: corrected=192;
219: corrected=193;
220: corrected=195;
221: corrected=197;
222: corrected=198;
223: corrected=200;
224: corrected=201;
225: corrected=203;
226: corrected=205;
227: corrected=206;
228: corrected=208;
229: corrected=210;
230: corrected=211;
231: corrected=213;
232: corrected=215;
233: corrected=216;
234: corrected=218;
235: corrected=220;
236: corrected=221;
237: corrected=223;
238: corrected=225;
239: corrected=226;
240: corrected=228;
241: corrected=230;
242: corrected=232;
243: corrected=233;
244: corrected=235;
245: corrected=237;
246: corrected=239;
247: corrected=240;
248: corrected=242;
249: corrected=244;
250: corrected=246;
251: corrected=247;
252: corrected=249;
253: corrected=251;
254: corrected=253;
255: corrected=255;


endcase 

endmodule

